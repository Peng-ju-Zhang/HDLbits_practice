`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/08/02 17:27:29
// Design Name: 
// Module Name: verilog
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module verilog_tb();
reg a,b,c;
wire w,x,y,z;
initial begin
a=0;b=1;c=0;
end
always #2 {a,b,c}={~a,~b,~c};

top_module top_module_tb(
	a,b,c
	,w,x,y,z);
endmodule